///////////////////////////////////////////////////////////////////////
// Write a 32-bit ripple-carry adder.
// 
// Implement your adder it by instantiating 32 1-bit full adders (fa1)
// and connecting them properly.  You can either instantiate them
// explicitely or as an array of modules or using generate statements.
//
// The signal names are self-explanatory.
///////////////////////////////////////////////////////////////////////

module FA32(a, b, cin, sum, cout);

  input  [31:0] a, b;
  input  cin;
  output [31:0] sum;
  output cout;
  
  
endmodule // top


